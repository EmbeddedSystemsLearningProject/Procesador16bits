module sumador (
    input  [7:0] inA,
    input  [7:0] inB,
    output [7:0] out
);

assign out = inA;
endmodule